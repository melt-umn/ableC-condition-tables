grammar edu:umn:cs:melt:exts:ableC:tables;

exports edu:umn:cs:melt:exts:ableC:tables:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:tables:abstractsyntax;

