grammar edu:umn:cs:melt:exts:ableC:tables:abstractsyntax;

imports edu:umn:cs:melt:ableC:abstractsyntax:host as abs;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction as abs;
imports edu:umn:cs:melt:ableC:abstractsyntax:env as abs;

imports silver:langutil;
imports silver:langutil:pp;

abstract production table
top::abs:Expr ::= trows::TableRows
{
  top.pp = ppConcat( [text("table ("), line(), trows.pp, text(" )")] );
  propagate abs:env, abs:controlStmtContext;

  forwards to 
    if !null(trows.errors) then
      abs:errorExpr(trows.errors, location=trows.location)
    else
      abs:stmtExpr(
        abs:foldStmt(trows.preDecls),
        disjunction(mapConjunction(transpose(trows.ftExprss))),
        location=top.location);
}

-- Table Rows --
----------------
nonterminal TableRows with pp, errors, abs:env, location,
  ftExprss, rlen, preDecls, abs:controlStmtContext;
propagate abs:env, abs:controlStmtContext on TableRows;

synthesized attribute preDecls :: [abs:Stmt];
synthesized attribute ftExprss :: [[abs:Expr]];
synthesized attribute rlen :: Integer;

abstract production tableRowSnoc
top::TableRows ::= trowstail::TableRows  trow::TableRow
{
  top.pp = ppConcat([trowstail.pp, line(), trow.pp]);

  top.errors := trowstail.errors ++ trow.errors;
  top.errors <-
    if trow.rlen == trowstail.rlen then [] else
      [err(trowstail.location,
        "The number of T,F,* entries in table row must be the same " ++
        "as the preceding rows")];

  top.rlen = trow.rlen;
  top.ftExprss = trowstail.ftExprss ++ [trow.ftExprs];
  top.preDecls = trowstail.preDecls ++ trow.preDecls;
}

abstract production tableRowOne
top::TableRows ::= trow::TableRow
{
  top.pp = trow.pp;
  top.errors := trow.errors;
  top.rlen = trow.rlen;
  top.ftExprss = [trow.ftExprs];
  top.preDecls = trow.preDecls;
}

-- Table Row --
---------------
nonterminal TableRow with pp, errors, abs:env, location,
  ftExprs, rlen, preDecls, abs:controlStmtContext;
propagate abs:env, abs:controlStmtContext on TableRow;

synthesized attribute ftExprs :: [abs:Expr];

abstract production tableRow
top::TableRow ::= e::abs:Expr tvl::TruthFlagList
{
  top.pp = ppConcat([e.pp, text(" : "), tvl.pp]);
  top.errors := e.errors;
  top.rlen = tvl.rlen;
  top.ftExprs = tvl.ftExprs;
  
  top.errors <-
    if abs:typeAssignableTo(abs:builtinType(abs:nilQualifier(), abs:boolType()), e.abs:typerep) then []
    else [err(e.location, "Condition expression expected type boolean (got " ++ abs:showType(e.abs:typerep) ++ ")")];
  
  -- Generate a name
  local ident :: abs:Name =
    abs:name("__table_condition_" ++ toString(genInt()), location = top.location);
  
  top.preDecls =
    [abs:declStmt(
      abs:variableDecls(
        abs:nilStorageClass(),
        abs:nilAttribute(),
        abs:directTypeExpr(
          abs:builtinType(abs:nilQualifier(), abs:boolType())),
        abs:foldDeclarator([
          abs:declarator(
            ident,
            abs:baseTypeExpr(),
            abs:nilAttribute(),
            abs:justInitializer(
              abs:exprInitializer(e, location=top.location))
          )
        ])
      )
    )]; -- _Bool ident = e;
  
  tvl.rowExpr = 
    abs:declRefExpr(ident, location=top.location);
}

-- Truth Value List
-------------------
nonterminal TruthFlagList with pp, rowExpr, ftExprs, rlen;

inherited attribute rowExpr :: abs:Expr;
-- the expression in the table row.  It is passed down to the TF*
-- values to be used in the translation to the host language.

abstract production tvlistCons
top::TruthFlagList ::= tv::TruthFlag  tvltail::TruthFlagList
{
  top.pp = ppConcat([tv.pp, text(" "), tvltail.pp]);
  top.rlen = 1 + tvltail.rlen;
  top.ftExprs = tv.ftExpr :: tvltail.ftExprs;

  tv.rowExpr = top.rowExpr;
  tvltail.rowExpr = top.rowExpr;
}

abstract production tvlistOne
top::TruthFlagList ::= tv::TruthFlag
{
  top.pp = tv.pp;
  top.rlen = 1;
  top.ftExprs = [tv.ftExpr];
 
  tv.rowExpr = top.rowExpr;
}


-- Truth Values
---------------
nonterminal TruthFlag with pp, rowExpr, ftExpr;

synthesized attribute ftExpr :: abs:Expr;

abstract production tvTrue
top::TruthFlag ::=
{
  top.pp = text("T");
  top.ftExpr = top.rowExpr;
}

abstract production tvFalse
top::TruthFlag ::=
{
  top.pp = text("F");
  top.ftExpr = logicalNegate(top.rowExpr);
}

abstract production tvStar
top::TruthFlag ::=
{ 
  top.pp = text("*");
  top.ftExpr =
    abs:realConstant(
      abs:integerConstant("1", false, abs:noIntSuffix(), location=top.rowExpr.location),
      location=top.rowExpr.location);
}


-- Our AST construction helper functions

function logicalNegate
abs:Expr ::= ne::abs:Expr
{
  return abs:notExpr(ne, location=ne.location);
}
function logicalOr
abs:Expr ::= e1::abs:Expr e2::abs:Expr
{
  return abs:orExpr(e1, e2, location=e1.location);
}
function logicalAnd
abs:Expr ::= e1::abs:Expr e2::abs:Expr
{
  return abs:andExpr(e1, e2, location=e1.location);
}

-- table helper functions
-------------------------
function disjunction
abs:Expr ::= es::[abs:Expr]
{
  return if length(es) == 1 then head(es)
         else logicalOr(head(es), disjunction(tail(es)));
}
function mapConjunction
[abs:Expr] ::= ess::[[abs:Expr]]
{
  return if null(ess) then [] 
         else cons(conjunction(head(ess)),
                     mapConjunction(tail(ess)));
}
function conjunction
abs:Expr ::= es::[abs:Expr]
{
  return if length(es) == 1 then head(es)
         else logicalAnd(head(es), conjunction(tail(es)));
}
function transpose
[[a]] ::= m::[[a]]
{
  return
    case m of
    | [] :: _ -> []
    | _       -> map(head,m) :: transpose(map(tail,m))
    end;
}

